library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

entity ROM is
    Port (
        clk       : in  std_logic;
        write     : in  std_logic;
        disable   : in  std_logic;
        address   : in  std_logic_vector(11 downto 0);
        datain    : in  std_logic_vector(35 downto 0);
        dataout   : out std_logic_vector(35 downto 0)
          );
end ROM; 

architecture Behavioral of ROM is

type memory_array is array (0 to ((2 ** 12) - 1) ) of std_logic_vector (35 downto 0); 

signal memory : memory_array:= (
--20 son opcodes & 16 son literales (o 12 son direcciones {11 downto 0})
	"000000000000000001000000000000000101",  -- MOV A,Lit(5)
	"000000000000000010000000000000000011",  -- MOV B,Lit(3)
	"000000000000000000110000000000000000",  -- MOV(Dir=0x00),B
	"000000000000010000110000000000000001",  -- SUB A,Lit(1)
	"000000000000010110000000000000000000",  -- CMP A,Lit(0)
	"000000000000010100000000000000001011",  -- JEQ (0x11)
	"000000000000010000000000000000000001",  -- MOV (Dir=0x01),A
	"000000000000000000010000000000000000",  -- MOV A,B
	"000000000000000001110000000000000000",  -- ADD B,(Dir=0x00)
	"000000000000000100000000000000000001",  -- MOV A,(Dir=0x01)
	"000000000000001100000000000000000011",  -- JMP (0x03)
	"000000000000000000000000000000000000",  -- NOP
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000",
	"000000000000000000000000000000000000"
        ); 

begin

process (clk)
    begin
       if (rising_edge(clk)) then
            if(write = '1') then
                memory(to_integer(unsigned(address))) <= datain;
            end if;
       end if;
end process;

with disable select
    dataout <= memory(to_integer(unsigned(address)))  when '0',
            (others => '0') when others;
            
end Behavioral; 

